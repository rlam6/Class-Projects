LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;

ENTITY mux21 IS
	GENERIC (NBIT : INTEGER := 32);
	PORT (	D1, D0 : IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
		S: IN STD_LOGIC;
		Y : OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0));
END ENTITY;

ARCHITECTURE mux21 OF mux21 IS
BEGIN
       Y <= D1 WHEN S='1' ELSE D0;
END ARCHITECTURE;
