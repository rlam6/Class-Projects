 --------------------------MUX DEFINITION----------------------------------------
LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX41 IS
	GENERIC(NBIT: INTEGER := 32);
	PORT(D3, D2, D1, D0 : IN STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0);
	     S   	    : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
	     Y              : OUT STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0));
END MUX41;

ARCHITECTURE MUX41 OF MUX41 IS
BEGIN
	Y <= D0 WHEN S = "00" ELSE
	     D1 WHEN S = "01" ELSE
	     D2 WHEN S = "10" ELSE
	     D3 WHEN S = "11";
END ARCHITECTURE;

LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
ENTITY MUX83 IS
	GENERIC(NBIT: INTEGER := 32);
	PORT(D7, D6, D5, D4, D3, D2, D1, D0: IN STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0);
	     S  		           : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	     Y  			   : OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0));
END MUX83;

ARCHITECTURE MUX83 OF MUX83 IS
COMPONENT MUX41 IS
	PORT(D3, D2, D1, D0 : IN STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0);
	     S   	    : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
	     Y              : OUT STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0));
END COMPONENT;
SIGNAL Y1, Y2 : STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0);
BEGIN
	Y1SEL : MUX41 PORT MAP (D7, D6, D5, D4, S(1 DOWNTO 0), Y1);
	Y2SEL : MUX41 PORT MAP (D3, D2, D1, D0, S(1 DOWNTO 0), Y2);
	Y <= Y1 WHEN S(2) = '1' ELSE Y2;
END ARCHITECTURE;

LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
ENTITY MUX81 IS
	PORT(D7, D6, D5, D4, D3, D2, D1, D0: IN STD_LOGIC;
	     S  		           : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	     Y  			   : OUT STD_LOGIC);
END MUX81;

ARCHITECTURE MUX81 OF MUX81 IS
BEGIN
	Y <= D0 WHEN S = "000" ELSE
	     D1 WHEN S = "001" ELSE
	     D2 WHEN S = "010" ELSE
	     D3 WHEN S = "011" ELSE
	     D4 WHEN S = "100" ELSE
	     D5 WHEN S = "101" ELSE
	     D6 WHEN S = "110" ELSE
	     D7 WHEN S = "111"; 
END ARCHITECTURE;
	
--------------------------Full-Adder (FA) Definition----------------------------
LIBRARY ieee;
	USE ieee.std_logic_1164.ALL;

ENTITY FA IS
	PORT(i0, i1, cin: IN STD_LOGIC; s, cout: OUT STD_LOGIC);
END FA;

ARCHITECTURE FA_Arch OF FA IS
BEGIN
	s <= (NOT i0 AND NOT i1 AND cin) OR
		(NOT i0 AND i1 AND NOT cin) OR
		(i0 AND NOt i1 AND NOT cin) OR
		(i0 AND i1 AND cin);
	
	cout <=	(NOT i0 AND i1 AND cin) OR
			(i0 AND NOT i1 AND cin) OR
			(i0 AND i1 AND NOT cin) OR
			(i0 AND i1 AND cin);
END FA_Arch;
-----------------COMPARATOR32-----------------------
LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;

ENTITY COMP32 IS
	GENERIC(NBIT : INTEGER := 32);
	PORT(A, B: IN STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0); 
	     GT, LT, EQ: OUT STD_LOGIC
		);
END ENTITY;
ARCHITECTURE COMP1 OF COMP32 IS
BEGIN
	GT <= '1' WHEN (A > B) ELSE '0';
	LT <= '1' WHEN (A < B) ELSE '0';
	EQ <= '1' WHEN (A = B) ELSE '0';
END ARCHITECTURE;
------------------------NOT 32--------------------------
LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;

ENTITY NOT32 IS
	GENERIC(NBIT: INTEGER := 32);
	PORT(A: IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0); 
	     Y: OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0)
		);
END NOT32;
ARCHITECTURE NOT_Arch OF NOT32 IS
BEGIN
	NOT4 : FOR I IN NBIT-1 DOWNTO 0 GENERATE
	BEGIN
		Y(I) <= NOT A(I);
	END GENERATE;
END ARCHITECTURE;
------------------------FA 32--------------------------
LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FA32 IS
	GENERIC(NBIT: INTEGER := 32);
	PORT(A, B: IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0); 
	     Y: OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	     COUT : OUT STD_LOGIC);
END FA32;
ARCHITECTURE FA_Arch OF FA32 IS
COMPONENT FA IS
	PORT(i0, i1, cin: IN STD_LOGIC; s, cout: OUT STD_LOGIC);
END COMPONENT;
SIGNAL CIN : STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0) := (OTHERS => '0');
BEGIN
	ADD31 : FOR I IN 0 TO NBIT-2 GENERATE
	BEGIN
		ADD : FA PORT MAP (A(I), B(I), CIN(I), Y(I), CIN(I+1));
	END GENERATE;
	LAST : FA PORT MAP (A(NBIT-1), B(NBIT-1), CIN(NBIT-1), Y(NBIT-1), COUT);
END ARCHITECTURE;

------------------------SUB4---------------------------
LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SUB32 IS
	GENERIC(NBIT: INTEGER := 32);
	PORT(A, B: IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0); 
	     Y: OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	     DOUT : OUT STD_LOGIC);
END ENTITY;
ARCHITECTURE SUB32 OF SUB32 IS
COMPONENT NOT32 IS
	PORT(A: IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0); Y: OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0));
END COMPONENT;
COMPONENT FA IS
	PORT(i0, i1, cin: IN STD_LOGIC; s, cout: OUT STD_LOGIC);
END COMPONENT;
SIGNAL DIN : STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0) := (0 => '1', OTHERS => '0');
SIGNAL BFIX : STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
BEGIN
	NOTB : NOT32 PORT MAP (B, BFIX);
	SUB31 : FOR I IN 0 TO NBIT-2 GENERATE
	BEGIN
		ADD : FA PORT MAP (A(I), BFIX(I), DIN(I), Y(I), DIN(I+1));
	END GENERATE;
	LAST : FA PORT MAP (A(NBIT-1), BFIX(NBIT-1), DIN(NBIT-1), Y(NBIT-1), DOUT);
END ARCHITECTURE;
------------------------SUBC4---------------------------
LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
ENTITY SUBC32 IS
	GENERIC(NBIT: INTEGER := 32);
	PORT(A, B: IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0); 
	     Y: OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	     DOUT : OUT STD_LOGIC);
END ENTITY;
ARCHITECTURE SUBC32 OF SUBC32 IS
COMPONENT NOT32 IS
	PORT(A: IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0); Y: OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0));
END COMPONENT;
COMPONENT FA IS
	PORT(i0, i1, cin: IN STD_LOGIC; s, cout: OUT STD_LOGIC);
END COMPONENT;
SIGNAL DIN : STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0) := (OTHERS => '0');
SIGNAL BFIX : STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
BEGIN
	NOTB : NOT32 PORT MAP (B, BFIX);
	SUBC31 : FOR I IN 0 TO NBIT-2 GENERATE
	BEGIN
		ADD : FA PORT MAP (A(I), BFIX(I), DIN(I), Y(I), DIN(I+1));
	END GENERATE;
	LAST : FA PORT MAP (A(NBIT-1), BFIX(NBIT-1), DIN(NBIT-1), Y(NBIT-1), DOUT);
END ARCHITECTURE;
------------------------MOVE32---------------------------
LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MOVE32 IS
	GENERIC(NBIT: INTEGER := 32);
	PORT(A: IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0); 
	     Y: OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0)
	);
END ENTITY;
ARCHITECTURE MOVE32 OF MOVE32 IS
BEGIN
	MOVE: FOR I IN NBIT-1 DOWNTO 0 GENERATE
	BEGIN
		Y(I) <= A(I);
	END GENERATE;
END ARCHITECTURE;
------------------------INC----------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY INC IS
	GENERIC(NBIT: INTEGER := 32);
	PORT (SIGNAL A : IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL Y : OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL COUT : OUT STD_LOGIC
		);
END ENTITY;
ARCHITECTURE INC OF INC IS
SIGNAL B : STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0) := (0 => '1', OTHERS => '0');
SIGNAL CIN : STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0) := (OTHERS => '0');
COMPONENT FA IS
	PORT(i0, i1, cin: IN STD_LOGIC; s, cout: OUT STD_LOGIC);
END COMPONENT;
BEGIN
	INCR : FOR i IN 0 TO NBIT-2 GENERATE
	BEGIN	
		ADD : FA PORT MAP (A(i), B(i), CIN(i), Y(i), CIN(i+1));
	END GENERATE;
	LAST : FA PORT MAP (A(NBIT-1), B(NBIT-1), CIN(NBIT-1), Y(NBIT-1), COUT);
END ARCHITECTURE;
------------------------DEC----------------------------
LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
ENTITY DEC32 IS
	GENERIC(NBIT: INTEGER := 32);
	PORT (SIGNAL A : IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL Y : OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL DOUT : OUT STD_LOGIC
		);
END ENTITY;
ARCHITECTURE DEC OF DEC32 IS
COMPONENT SUB32 IS
	PORT(A, B: IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0); Y: OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	     DOUT : OUT STD_LOGIC);
END COMPONENT;
SIGNAL B : STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0) := (0 => '1', OTHERS => '0');
BEGIN
	DECR : SUB32 PORT MAP (A, B, Y, DOUT);
END ARCHITECTURE;
------------------------ADDINC----------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY ADDINC IS
	GENERIC(NBIT: INTEGER := 32);
	PORT (SIGNAL A, B : IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL Y : OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL COUT : OUT STD_LOGIC
		);
END ENTITY;
ARCHITECTURE ADDINC OF ADDINC IS
SIGNAL CIN1, CIN2 : STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0) := (OTHERS => '0');
SIGNAL Y1 : STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
SIGNAL CEXTRA : STD_LOGIC;
COMPONENT FA32 IS
	PORT(A, B: IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0); 
	     Y: OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	     COUT : OUT STD_LOGIC);
END COMPONENT;
COMPONENT INC IS
	PORT (SIGNAL A : IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL Y : OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL COUT : OUT STD_LOGIC
		);
END COMPONENT;
BEGIN
	ADD : FA32 PORT MAP (A, B, Y1, CEXTRA);
	INCR : INC PORT MAP (Y1, Y, COUT);
END ARCHITECTURE;
------------------------AND--------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY ANDGATE IS
	GENERIC(NBIT: INTEGER := 32);
	PORT (SIGNAL A, B : IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL Y : OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0)
		);
END ENTITY;
ARCHITECTURE ANDGATE OF ANDGATE IS
BEGIN
	ANDRUN : FOR I IN NBIT-1 DOWNTO 0 GENERATE
	BEGIN
		Y(I) <= A(I) AND B(I);
	END GENERATE;
END ARCHITECTURE;
------------------------OR--------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY ORGATE IS
	GENERIC(NBIT: INTEGER := 32);
	PORT (SIGNAL A, B : IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL Y : OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0)
		);
END ENTITY;
ARCHITECTURE ORGATE OF ORGATE IS
BEGIN
	ORRUN : FOR I IN NBIT-1 DOWNTO 0 GENERATE
	BEGIN
		Y(I) <= A(I) OR B(I);
	END GENERATE;
END ARCHITECTURE;
------------------------XOR--------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY XORGATE IS
	GENERIC(NBIT: INTEGER := 32);
	PORT (SIGNAL A, B : IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL Y : OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0)
		);
END ENTITY;
ARCHITECTURE XORGATE OF XORGATE IS
BEGIN
	XORRUN : FOR I IN NBIT-1 DOWNTO 0 GENERATE
	BEGIN
		Y(I) <= A(I) XOR B(I);
	END GENERATE;
END ARCHITECTURE;
------------------------SHL--------------------------------
LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
	USE IEEE.NUMERIC_STD.ALL;
ENTITY SHL IS
	GENERIC(NBIT: INTEGER := 32; STEP : INTEGER := 1);
	PORT (SIGNAL A, B : IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL Y    : OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0)
		);
END ENTITY;
ARCHITECTURE SHL OF SHL IS
BEGIN
	SHIFT : FOR I IN NBIT-STEP-1 DOWNTO 0 GENERATE
	BEGIN
		Y(I+STEP) <= A(I);
	END GENERATE;
	ADD_ZEROS : FOR I IN STEP-1 DOWNTO 0 GENERATE
	BEGIN
		Y(I) <= '0';
	END GENERATE;
END ARCHITECTURE;
------------------------COMP--------------------------------
LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
ENTITY COMP IS
	GENERIC(NBIT: INTEGER := 32);
	PORT (SIGNAL A, B : IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL Y    : OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0)
		);
END ENTITY;
ARCHITECTURE COMP OF COMP IS
BEGIN
	COMPARE : FOR I IN NBIT-1 DOWNTO 0 GENERATE
	BEGIN
		Y(I) <= '1' WHEN (A(I) > B(I)) ELSE '0';
	END GENERATE;
END ARCHITECTURE;
------------------------ALU--------------------------------
LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
	USE IEEE.STD_LOGIC_ARITH.ALL;
	USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY ALU IS
	GENERIC(NBIT: INTEGER := 32);
	PORT (SIGNAL A, B : IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL R    : IN STD_LOGIC;
	      SIGNAL FUNCT : STD_LOGIC_VECTOR (3 DOWNTO 0);
	      SIGNAL OUTPUT : OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL COUT, EQUAL, OVERFLOW : OUT STD_LOGIC
		);
END ENTITY;
ARCHITECTURE ALU OF ALU IS
COMPONENT MUX81 IS
	PORT(D7, D6, D5, D4, D3, D2, D1, D0 : IN STD_LOGIC;
	     S   : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
	     Y   : OUT STD_LOGIC);
END COMPONENT;
COMPONENT MUX83 IS
	PORT(D7, D6, D5, D4, D3, D2, D1, D0 : IN STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0);
	     S   : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
	     Y   : OUT STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0));
END COMPONENT;
COMPONENT COMP32 IS
	PORT(A, B: IN STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0); 
	     GT, LT, EQ: OUT STD_LOGIC
		);
END COMPONENT;
COMPONENT NOT32 IS
	PORT(A: IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0); 
	     Y: OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0)
		);
END COMPONENT;
COMPONENT FA32 IS
	PORT(A, B: IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0); 
	     Y: OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	     COUT : OUT STD_LOGIC);
END COMPONENT;
COMPONENT SUB32 IS
	PORT(A, B: IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0); 
	     Y: OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	     DOUT : OUT STD_LOGIC);
END COMPONENT;
COMPONENT SUBC32 IS
	PORT(A, B: IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0); 
	     Y: OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	     DOUT : OUT STD_LOGIC);
END COMPONENT;
COMPONENT MOVE32 IS
	PORT(A: IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0); 
	     Y: OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0));
END COMPONENT;
COMPONENT INC IS
	PORT (SIGNAL A : IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL Y : OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL COUT : OUT STD_LOGIC
		);
END COMPONENT;
COMPONENT DEC32 IS
	PORT (SIGNAL A : IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL Y : OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL DOUT : OUT STD_LOGIC);
END COMPONENT;
COMPONENT ADDINC IS
	PORT (SIGNAL A, B : IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL Y : OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL COUT : OUT STD_LOGIC);
END COMPONENT;
COMPONENT ANDGATE IS
	PORT (SIGNAL A, B : IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL Y : OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0)
		);
END COMPONENT;
COMPONENT ORGATE IS
	PORT (SIGNAL A, B : IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL Y : OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0)
		);
END COMPONENT;
COMPONENT XORGATE IS
	PORT (SIGNAL A, B : IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL Y : OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0)
		);
END COMPONENT;
COMPONENT SHL IS
	GENERIC(NBIT: INTEGER := 32; STEP : INTEGER := 1);
	PORT (SIGNAL A, B : IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL Y : OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0)
		);
END COMPONENT;
COMPONENT COMP IS
	GENERIC(NBIT: INTEGER := 32);
	PORT (SIGNAL A, B : IN STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
	      SIGNAL Y    : OUT STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0)
		);
END COMPONENT;
---------------------BEGIN SIGNAL DECLARATIONS----------------------
SIGNAL addComp, subcComp, move0, move1, move, subComp : STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
SIGNAL incComp, decComp, addincrComp, compareComp : STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
SIGNAL andComp, orComp, xorComp, complComp, bitSHLComp : STD_LOGIC_VECTOR (NBIT-1 DOWNTO 0);
SIGNAL addCOUT, subcCOUT, incCOUT, decCOUT, addincrCOUT : STD_LOGIC;
SIGNAL bitSHLCOUT, subCOUT, dontCareOne, cout0, cout1 : STD_LOGIC;
SIGNAL dontCare, sel1, sel0: STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0);
SIGNAL greaterthan, lessthan : STD_LOGIC;
SIGNAL MODE : STD_LOGIC;
SIGNAL opsel : STD_LOGIC_VECTOR (2 DOWNTO 0);
---------------------END SIGNAL DECLARATIONS------------------------
BEGIN
	MODE <= FUNCT(3); opsel <= FUNCT(2 DOWNTO 0);
	dontCare <= (OTHERS => 'X');
	dontCareOne <= 'X';
	-------------SELECT PORT INPUTS--------------------
	add      : FA32 PORT MAP (A, B, addComp, addCOUT);
	subBC    : SUBC32 PORT MAP (A, B, subcComp, subcCOUT);
	subtract : SUB32 PORT MAP (A, B, subComp, subCOUT);
	incr     : INC PORT MAP (A, incComp, incCOUT);
	decr     : DEC32 PORT MAP (A, decComp, decCOUT);
	addincr  : ADDINC PORT MAP (A, B, addincrComp, addincrCOUT);
	orG      : ORGATE PORT MAP (A, B, orComp);
	andG     : ANDGATE PORT MAP (A, B, andComp);
	xorG     : XORGATE PORT MAP (A, B, xorComp);
	move0Comp: MOVE32 PORT MAP (A, move0);
	move1Comp: MOVE32 PORT MAP (B, move1);
	compG    : NOT32 PORT MAP (A, complComp);
	BITSHL   : SHL PORT MAP (A, B, bitSHLComp);
	compareG : COMP PORT MAP (A, B, compareComp);
	compaG   : COMP32 PORT MAP (A, B, greaterthan, lessthan, EQUAL);

	move <= move0 WHEN R='1' ELSE move1;
	-------------OUTPUTS SELECTIONS----------------------------------
	MUX81A : MUX83 PORT MAP (complComp, orComp, andComp, dontCare, compareComp,
				subComp, addComp, dontCare, opsel, sel0);
	MUX81B : MUX83 PORT MAP (dontCare, dontCare, dontCare, dontCare, move,
				dontCare, bitSHLComp, xorComp, opsel, sel1);

	-------------COUT SELECTIONS--------------------------------------
	MUX81C : MUX81 PORT MAP (dontCareOne, dontCareOne, dontCareOne, dontCareOne,
				dontCareOne, subCOUT, addCOUT, dontCareOne,
				opsel, cout0);
	MUX81D : MUX81 PORT MAP (dontCareOne, dontCareOne, dontCareOne, dontCareOne,
				dontCareOne, dontCareOne, bitSHLCOUT, dontCareOne,
				opsel, cout1);
	-------------OUTPUTS---------------------
	OUTPUT   <= sel1 WHEN MODE='1' ELSE sel0;
	COUT     <= cout1 WHEN MODE='1' ELSE cout0;
	OVERFLOW <= '1' WHEN (cout1 = '1' OR cout0 = '1') ELSE '0';

END ARCHITECTURE;
